//Verilog HDL for ""0814_opamp_N_P, ""
`timescale 1 ps / 1 ps

module X0814_opamp_N_P ( 
  inout wire VOUT,
  input wire VINm, VINp 
  );

//   pullup (weak1) pu1 (REF);
//   pullup (weak1) pu1 (FRCREF);
   

endmodule
