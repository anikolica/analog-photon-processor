VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO pathCL STRING ;
  MACRO arrayDisplay STRING ;
  MACRO instLabel STRING ;
  MACRO startLevel INTEGER ;
  MACRO stopLevel INTEGER ;
  MACRO scrollPercent INTEGER ;
  MACRO gridSpacing REAL ;
  MACRO gridMultiple INTEGER ;
  MACRO xSnapSpacing REAL ;
  MACRO ySnapSpacing REAL ;
  MACRO snapMode STRING ;
  MACRO segSnapMode STRING ;
  MACRO instanceDrawingMode STRING ;
  MACRO lppVisibilityMode STRING ;
  MACRO filterSize REAL ;
  MACRO filterSizeDrawingStyle STRING ;
  MACRO displayResolution STRING ;
  MACRO dimmingScope STRING ;
  MACRO dimmingIntensity INTEGER ;
  MACRO autoZoomMode STRING ;
  MACRO autoZoomScale INTEGER ;
  MACRO mergeScope STRING ;
  MACRO viewNameList STRING ;
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER PDK
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.47 ;
  SPACING 0 LAYER NW ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.47 ;" ;
END PDK

LAYER NW
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_SPACING "SPACING 0.47 ;
  SPACING 2.5 LAYER DNW ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.47 ;" ;
END NW

LAYER OD
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE DIFFUSION ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.08 ;" ;
END OD

LAYER OD_33
  TYPE MASTERSLICE ;
END OD_33

LAYER OD_18
  TYPE MASTERSLICE ;
END OD_18

LAYER OD_25
  TYPE MASTERSLICE ;
END OD_25

LAYER PO
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.06 ;
  AREA 0.042 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 0.184 
    WIDTH 0.004 0.12 0.12 
    WIDTH 0.134 0.12 0.18 ;
  SPACING 0.12 SAMENET ;
  MINSTEP 0.08 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.094 ;
  DIAGSPACING 0.19 ;
  SPACING 0.14 ENDOFLINE 0.09 WITHIN 0.035 PARALLELEDGE 0.14 WITHIN 0.09 ;
  RESISTANCE RPERSQ 15.0619 ;
  CAPACITANCE CPERSQDIST 0.00637 ;
  THICKNESS 1000 ;
  EDGECAPACITANCE 0.0117 ;
  MINIMUMDENSITY 14 ;
  MAXIMUMDENSITY 40 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 250 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 250 ;
    ANTENNACUMAREARATIO 1000 ;
  PROPERTY LEF58_TYPE "TYPE POLYROUTING ;" ;
END PO

LAYER PP
  TYPE IMPLANT ;
  WIDTH 0.18 ;
  SPACING 0.18 ;
  AREA 0.122 ;
END PP

LAYER NP
  TYPE IMPLANT ;
  WIDTH 0.18 ;
  SPACING 0.18 ;
  AREA 0.122 ;
END NP

LAYER CO
  TYPE CUT ;
  SPACING 0.11 ;
  SPACING 0.14 ADJACENTCUTS 3 WITHIN 0.15 ;
  WIDTH 0.09 ;
  ENCLOSURE BELOW 0.01 0.04 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE ABOVE 0.04 0.04 WIDTH 1.005 ;
  ENCLOSURE ABOVE 0.025 0.025 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 10 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 10 ;
  PROPERTY LEF58_SPACING "SPACING 0.14 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END CO

LAYER M1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.18 0.18 ;
  WIDTH 0.09 ;
  OFFSET 0.09 0.09 ;
  AREA 0.042 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.419 1.499 4.499 
    WIDTH 0 0.09 0.09 0.09 0.09 0.09 
    WIDTH 0.2 0.09 0.11 0.11 0.11 0.11 
    WIDTH 0.42 0.09 0.11 0.16 0.16 0.16 
    WIDTH 1.5 0.09 0.11 0.16 0.5 0.5 
    WIDTH 4.5 0.09 0.11 0.16 0.5 1.5 ;
  SPACING 0.09 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.09 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.11 ENDOFLINE 0.11 WITHIN 0.035 PARALLELEDGE 0.11 WITHIN 0.11 ;
  RESISTANCE RPERSQ 0.0868 ;
  CAPACITANCE CPERSQDIST 0.00514 ;
  THICKNESS 1800 ;
  EDGECAPACITANCE 0.00758 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       9.36775 19.5501 39.9148 80.6441 253.744 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       1.20706 2.15515 3.93091 7.39472 21.9815 ;
END M1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  WIDTH 0.1 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE BELOW 0 0.04 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
  PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END VIA1

LAYER M2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.399 1.499 4.499 
    WIDTH 0 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.2 0.1 0.12 0.12 0.12 0.12 
    WIDTH 0.4 0.1 0.12 0.16 0.16 0.16 
    WIDTH 1.5 0.1 0.12 0.16 0.5 0.5 
    WIDTH 4.5 0.1 0.12 0.16 0.5 1.5 ;
  SPACING 0.1 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.1 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.00298 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00659 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.749923 1.31913 2.37142 4.41089 12.9754 ;
END M2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  WIDTH 0.1 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE BELOW 0 0.04 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
  PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END VIA2

LAYER M3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.399 1.499 4.499 
    WIDTH 0 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.2 0.1 0.12 0.12 0.12 0.12 
    WIDTH 0.4 0.1 0.12 0.16 0.16 0.16 
    WIDTH 1.5 0.1 0.12 0.16 0.5 0.5 
    WIDTH 4.5 0.1 0.12 0.16 0.5 1.5 ;
  SPACING 0.1 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.1 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.00199 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00578 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.696634 1.16947 1.99669 3.54867 9.95791 ;
END M3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  WIDTH 0.1 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE BELOW 0 0.04 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
  PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END VIA3

LAYER M4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.399 1.499 4.499 
    WIDTH 0 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.2 0.1 0.12 0.12 0.12 0.12 
    WIDTH 0.4 0.1 0.12 0.16 0.16 0.16 
    WIDTH 1.5 0.1 0.12 0.16 0.5 0.5 
    WIDTH 4.5 0.1 0.12 0.16 0.5 1.5 ;
  SPACING 0.1 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.1 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.00149 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00537 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.674844 1.10631 1.83204 3.15479 8.51792 ;
END M4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  WIDTH 0.1 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE BELOW 0 0.04 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
  PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END VIA4

LAYER M5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.399 1.499 4.499 
    WIDTH 0 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.2 0.1 0.12 0.12 0.12 0.12 
    WIDTH 0.4 0.1 0.12 0.16 0.16 0.16 
    WIDTH 1.5 0.1 0.12 0.16 0.5 0.5 
    WIDTH 4.5 0.1 0.12 0.16 0.5 1.5 ;
  SPACING 0.1 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.1 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.0012 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00513 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.59004 0.967284 1.60182 2.75834 7.44752 ;
END M5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  WIDTH 0.1 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE BELOW 0 0.04 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
  PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END VIA5

LAYER M6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.399 1.499 4.499 
    WIDTH 0 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.2 0.1 0.12 0.12 0.12 0.12 
    WIDTH 0.4 0.1 0.12 0.16 0.16 0.16 
    WIDTH 1.5 0.1 0.12 0.16 0.5 0.5 
    WIDTH 4.5 0.1 0.12 0.16 0.5 1.5 ;
  SPACING 0.1 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMABOVE LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMABOVE LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.1 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.000996 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00502 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.531302 0.870991 1.44236 2.48375 6.70612 ;
END M6

LAYER VIA6
  TYPE CUT ;
  SPACING 0.1 ;
  SPACING 0.13 ADJACENTCUTS 3 WITHIN 0.14 ;
  WIDTH 0.1 ;
  ENCLOSURE BELOW 0.03 0.03 ;
  ENCLOSURE BELOW 0 0.04 ;
  ENCLOSURE ABOVE 0.03 0.03 ;
  ENCLOSURE ABOVE 0 0.04 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
  PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ;" ;
END VIA6

LAYER M7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.2 0.2 ;
  WIDTH 0.1 ;
  OFFSET 0.1 0.1 ;
  AREA 0.052 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.379 0.399 1.499 4.499 
    WIDTH 0 0.1 0.1 0.1 0.1 0.1 
    WIDTH 0.2 0.1 0.12 0.12 0.12 0.12 
    WIDTH 0.4 0.1 0.12 0.16 0.16 0.16 
    WIDTH 1.5 0.1 0.12 0.16 0.5 0.5 
    WIDTH 4.5 0.1 0.12 0.16 0.5 1.5 ;
  SPACING 0.1 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 1.7 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.799 WITHIN 1.7 FROMABOVE ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 0.699 WITHIN 0.2 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.2 ;
  MINIMUMCUT 4 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.25 ;
  MINIMUMCUT 4 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.2 ;
  MINIMUMCUT 9 WIDTH 0.7 FROMBELOW LENGTH 0.7 WITHIN 0.35 ;
  MINIMUMCUT 2 WIDTH 0.3 FROMBELOW LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 2 WITHIN 2 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 1.8 FROMABOVE LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINSTEP 0.1 MAXEDGES 1 ;
  MINENCLOSEDAREA 0.2 ;
  DIAGPITCH 0.38 0.38 ;
  DIAGSPACING 0.19 ;
  SPACING 0.12 ENDOFLINE 0.12 WITHIN 0.035 PARALLELEDGE 0.12 WITHIN 0.12 ;
  RESISTANCE RPERSQ 0.0778 ;
  CAPACITANCE CPERSQDIST 0.000854 ;
  THICKNESS 2200 ;
  EDGECAPACITANCE 0.00529 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       5.72474 11.9473 24.3923 49.2825 155.066 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       0.486946 0.798276 1.32194 2.2764 6.14627 ;
END M7

LAYER VIA7
  TYPE CUT ;
  SPACING 0.34 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.02 0.08 ;
  ENCLOSURE ABOVE 0.02 0.08 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA7

LAYER M8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.8 0.8 ;
  WIDTH 0.4 ;
  OFFSET 0.4 0.4 ;
  AREA 0.565 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0.004 1.504 4.504 
    WIDTH 0.004 0.4 0.4 0.4 
    WIDTH 1.504 0.4 0.5 0.5 
    WIDTH 4.504 0.4 0.5 1.5 ;
  SPACING 0.4 SAMENET ;
  MINIMUMCUT 1 WIDTH 0 WITHIN 1.7 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.799 WITHIN 1.7 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0 WITHIN 1.7 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.8 FROMBELOW LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 1.8 FROMABOVE LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMABOVE LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 0.565 ;
  RESISTANCE RPERSQ 0.0215 ;
  CAPACITANCE CPERSQDIST 0.00323 ;
  THICKNESS 9000 ;
  EDGECAPACITANCE 0.00615 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 90 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       16.0372 33.8563 69.4945 140.771 443.695 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       1.29043 2.05444 3.2317 5.20772 12.6666 ;
END M8

LAYER VIA8
  TYPE CUT ;
  SPACING 0.34 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.56 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.08 0.08 ;
  ENCLOSURE ABOVE 0.3 0.3 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 20 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNAAREARATIO 20 ;
END VIA8

LAYER M9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 4 4 ;
  WIDTH 2 ;
  OFFSET 2 2 ;
  AREA 9 ;
  SPACING 2 ;
  SPACING 2 SAMENET ;
  MINIMUMCUT 2 WIDTH 0 WITHIN 1.7 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.8 FROMBELOW LENGTH 1.8 WITHIN 1.7 ;
  MINIMUMCUT 2 WIDTH 3 FROMBELOW LENGTH 10 WITHIN 5 ;
  MAXWIDTH 12 ;
  MINENCLOSEDAREA 9 ;
  RESISTANCE RPERSQ 0.0215 ;
  CAPACITANCE CPERSQDIST 0.00245 ;
  THICKNESS 34000 ;
  EDGECAPACITANCE 0.00564 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 80 ;
  DENSITYCHECKWINDOW 75 75 ;
  DENSITYCHECKSTEP 37.5 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
  ACCURRENTDENSITY PEAK
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       16.0372 33.8563 69.4945 140.771 443.695 ;
  ACCURRENTDENSITY RMS
    FREQUENCY 1 ;
    WIDTH 0.2 0.4 0.8 1.6 5 ;
    TABLEENTRIES
       1.64281 2.60223 4.05931 6.46339 15.3636 ;
END M9

LAYER RV
  TYPE CUT ;
  SPACING 3 ;
  WIDTH 3 ;
  ENCLOSURE BELOW 1.5 1.5 ;
  ENCLOSURE ABOVE 1.5 1.5 ;
END RV

LAYER AP
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  WIDTH 3 ;
  SPACING 2 ;
  MAXWIDTH 35 ;
  MINIMUMDENSITY 10 ;
  MAXIMUMDENSITY 70 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNACUMAREARATIO 5000 ;
  ANTENNAMODEL OXIDE2 ;
    ANTENNACUMAREARATIO 1000 ;
END AP

MAXVIASTACK 4 RANGE M1 M7 ;
VIARULE AP_M9 GENERATE
  LAYER M9 ;
    ENCLOSURE 1.5 1.5 ;
  LAYER AP ;
    ENCLOSURE 1.5 1.5 ;
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
    SPACING 6 BY 6 ;
END AP_M9

VIARULE M9_M8 GENERATE DEFAULT
  LAYER M8 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER M9 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER VIA8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.7 BY 0.7 ;
END M9_M8

VIARULE M8_M7 GENERATE DEFAULT
  LAYER M7 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER M8 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.7 BY 0.7 ;
END M8_M7

VIARULE M7_M6 GENERATE DEFAULT
  LAYER M6 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M7 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M7_M6

VIARULE M6_M5 GENERATE DEFAULT
  LAYER M5 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M6 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M6_M5

VIARULE M5_M4 GENERATE DEFAULT
  LAYER M4 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M5 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M5_M4

VIARULE M4_M3 GENERATE DEFAULT
  LAYER M3 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M4 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M4_M3

VIARULE M3_M2 GENERATE DEFAULT
  LAYER M2 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M3 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M3_M2

VIARULE M2_M1 GENERATE DEFAULT
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M2 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
    SPACING 0.2 BY 0.2 ;
END M2_M1

VIARULE M1_PO GENERATE DEFAULT
  LAYER PO ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_PO

VIARULE M1_NPO GENERATE
  LAYER PO ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_NPO

VIARULE M1_PPO GENERATE
  LAYER PO ;
    ENCLOSURE 0.04 0.04 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_PPO

VIARULE M1_OD GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_OD

VIARULE M1_NOD GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_NOD

VIARULE M1_POD GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_POD

VIARULE M1_NW GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_NW

VIARULE M1_SUB GENERATE
  LAYER OD ;
    ENCLOSURE 0.03 0.03 ;
  LAYER M1 ;
    ENCLOSURE 0.04 0.04 ;
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
    SPACING 0.2 BY 0.2 ;
END M1_SUB

VIA DFM_M7_M6s
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M6 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M7_M6s

VIA DFM_M6_M5s
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M5 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M6_M5s

VIA DFM_M5_M4s
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M4 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M5_M4s

VIA DFM_M4_M3s
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M3 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M4_M3s

VIA DFM_M3_M2s
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M2 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M3_M2s

VIA DFM_M2_M1s
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.12 -0.12 0.12 0.12 ;
  LAYER M1 ;
    RECT -0.12 -0.12 0.12 0.12 ;
END DFM_M2_M1s

VIA DFM_M1_ODs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.105 -0.105 0.105 0.105 ;
  LAYER OD ;
    RECT -0.085 -0.085 0.085 0.085 ;
END DFM_M1_ODs

VIA DFM_M1_POs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.105 -0.105 0.105 0.105 ;
  LAYER PO ;
    RECT -0.105 -0.105 0.105 0.105 ;
END DFM_M1_POs

VIA AP_M9s
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER AP ;
    RECT -3 -3 3 3 ;
  LAYER M9 ;
    RECT -3 -3 3 3 ;
END AP_M9s

VIA M9_M8s
  LAYER VIA8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M9 ;
    RECT -0.58 -0.58 0.58 0.58 ;
  LAYER M8 ;
    RECT -0.26 -0.26 0.26 0.26 ;
END M9_M8s

VIA M8_M7s
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M8 ;
    RECT -0.26 -0.26 0.26 0.26 ;
  LAYER M7 ;
    RECT -0.26 -0.26 0.26 0.26 ;
END M8_M7s

VIA M7_M6s
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M7 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M6 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M7_M6s

VIA M6_M5s
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M5 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M6_M5s

VIA M5_M4s
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M4 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M5_M4s

VIA M4_M3s
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M3 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M4_M3s

VIA M3_M2s
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M2 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M3_M2s

VIA M2_M1s
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.09 -0.09 0.09 0.09 ;
  LAYER M1 ;
    RECT -0.09 -0.09 0.09 0.09 ;
END M2_M1s

VIA M1_ODs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER OD ;
    RECT -0.075 -0.075 0.075 0.075 ;
END M1_ODs

VIA M1_POs
  LAYER CO ;
    RECT -0.045 -0.045 0.045 0.045 ;
  LAYER M1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER PO ;
    RECT -0.085 -0.085 0.085 0.085 ;
END M1_POs

VIA M2_M1c
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M2 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M2_M1c

VIA M3_M2c
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M3 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M3_M2c

VIA M4_M3c
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M4 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M4_M3c

VIA M5_M4c
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M5 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M5_M4c

VIA M6_M5c
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M6 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M6_M5c

VIA M7_M6c
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.05 -0.09 0.05 0.09 ;
  LAYER M7 ;
    RECT -0.09 -0.05 0.09 0.05 ;
END M7_M6c

VIA M8_M7c
  LAYER VIA7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M7 ;
    RECT -0.2 -0.26 0.2 0.26 ;
  LAYER M8 ;
    RECT -0.26 -0.2 0.26 0.2 ;
END M8_M7c

VIA M9_M8c
  LAYER VIA8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER M8 ;
    RECT -0.48 -0.26 0.48 0.26 ;
  LAYER M9 ;
    RECT -0.26 -0.48 0.26 0.48 ;
END M9_M8c

VIA AP_M9c
  LAYER RV ;
    RECT -1.5 -1.5 1.5 1.5 ;
  LAYER M9 ;
    RECT -3 -3 3 3 ;
  LAYER AP ;
    RECT -3 -3 3 3 ;
END AP_M9c

VIA DFM_M2_M1c
  LAYER VIA1 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M1 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M2 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M2_M1c

VIA DFM_M3_M2c
  LAYER VIA2 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M2 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M3 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M3_M2c

VIA DFM_M4_M3c
  LAYER VIA3 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M3 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M4 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M4_M3c

VIA DFM_M5_M4c
  LAYER VIA4 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M4 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M5 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M5_M4c

VIA DFM_M6_M5c
  LAYER VIA5 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M5 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M6 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M6_M5c

VIA DFM_M7_M6c
  LAYER VIA6 ;
    RECT -0.05 -0.05 0.05 0.05 ;
  LAYER M6 ;
    RECT -0.09 -0.12 0.09 0.12 ;
  LAYER M7 ;
    RECT -0.12 -0.09 0.12 0.09 ;
END DFM_M7_M6c

NONDEFAULTRULE virtuosoDefaultSetup
  LAYER AP
    WIDTH 3 ;
  END AP
  LAYER M9
    WIDTH 2 ;
  END M9
  LAYER M8
    WIDTH 0.4 ;
  END M8
  LAYER M7
    WIDTH 0.1 ;
  END M7
  LAYER M6
    WIDTH 0.1 ;
  END M6
  LAYER M5
    WIDTH 0.1 ;
  END M5
  LAYER M4
    WIDTH 0.1 ;
  END M4
  LAYER M3
    WIDTH 0.1 ;
  END M3
  LAYER M2
    WIDTH 0.1 ;
  END M2
  LAYER M1
    WIDTH 0.09 ;
  END M1
  LAYER PO
    WIDTH 0.06 ;
  END PO
  USEVIARULE AP_M9 ;
  USEVIARULE M9_M8 ;
  USEVIARULE M8_M7 ;
  USEVIARULE M7_M6 ;
  USEVIARULE M6_M5 ;
  USEVIARULE M5_M4 ;
  USEVIARULE M4_M3 ;
  USEVIARULE M3_M2 ;
  USEVIARULE M2_M1 ;
  USEVIARULE M1_PO ;
  USEVIARULE M1_OD ;
  USEVIARULE M1_NPO ;
  USEVIARULE M1_PPO ;
  USEVIARULE M1_POD ;
  USEVIARULE M1_NOD ;
  USEVIARULE M1_NW ;
  USEVIARULE M1_SUB ;
END virtuosoDefaultSetup
NONDEFAULTRULE LEFDefaultRouteSpec_DFM
  LAYER M9
    WIDTH 2 ;
  END M9
  LAYER M8
    WIDTH 0.4 ;
  END M8
  LAYER M7
    WIDTH 0.1 ;
  END M7
  LAYER M6
    WIDTH 0.1 ;
  END M6
  LAYER M5
    WIDTH 0.1 ;
  END M5
  LAYER M4
    WIDTH 0.1 ;
  END M4
  LAYER M3
    WIDTH 0.1 ;
  END M3
  LAYER M2
    WIDTH 0.1 ;
  END M2
  LAYER M1
    WIDTH 0.09 ;
  END M1
  LAYER PO
    WIDTH 0.06 ;
  END PO
  USEVIARULE M9_M8 ;
  USEVIARULE M8_M7 ;
  USEVIARULE M7_M6 ;
  USEVIARULE M6_M5 ;
  USEVIARULE M5_M4 ;
  USEVIARULE M4_M3 ;
  USEVIARULE M3_M2 ;
  USEVIARULE M2_M1 ;
  USEVIARULE M1_PO ;
END LEFDefaultRouteSpec_DFM
MACRO X0814_opamp_N_P
  CLASS BLOCK ;
  ORIGIN 25.03 16.63 ;
  FOREIGN X0814_opamp_N_P -25.03 -16.63 ;
  SIZE 60 BY 65.005 ;
  SYMMETRY X Y R90 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 30.81 11.98 32.66 13.84 ;
      LAYER VIA2 ;
        RECT 30.72 13.7 30.82 13.8 ;
        RECT 30.72 13.46 30.82 13.56 ;
        RECT 30.72 13.22 30.82 13.32 ;
        RECT 30.72 12.98 30.82 13.08 ;
        RECT 30.72 12.74 30.82 12.84 ;
        RECT 30.72 12.5 30.82 12.6 ;
        RECT 30.72 12.26 30.82 12.36 ;
        RECT 30.72 12.02 30.82 12.12 ;
        RECT 30.92 13.7 31.02 13.8 ;
        RECT 30.92 13.46 31.02 13.56 ;
        RECT 30.92 13.22 31.02 13.32 ;
        RECT 30.92 12.98 31.02 13.08 ;
        RECT 30.92 12.74 31.02 12.84 ;
        RECT 30.92 12.5 31.02 12.6 ;
        RECT 30.92 12.26 31.02 12.36 ;
        RECT 30.92 12.02 31.02 12.12 ;
        RECT 31.12 13.7 31.22 13.8 ;
        RECT 31.12 13.46 31.22 13.56 ;
        RECT 31.12 13.22 31.22 13.32 ;
        RECT 31.12 12.98 31.22 13.08 ;
        RECT 31.12 12.74 31.22 12.84 ;
        RECT 31.12 12.5 31.22 12.6 ;
        RECT 31.12 12.26 31.22 12.36 ;
        RECT 31.12 12.02 31.22 12.12 ;
        RECT 31.32 13.7 31.42 13.8 ;
        RECT 31.32 13.46 31.42 13.56 ;
        RECT 31.32 13.22 31.42 13.32 ;
        RECT 31.32 12.98 31.42 13.08 ;
        RECT 31.32 12.74 31.42 12.84 ;
        RECT 31.32 12.5 31.42 12.6 ;
        RECT 31.32 12.26 31.42 12.36 ;
        RECT 31.32 12.02 31.42 12.12 ;
        RECT 31.52 13.7 31.62 13.8 ;
        RECT 31.52 13.46 31.62 13.56 ;
        RECT 31.52 13.22 31.62 13.32 ;
        RECT 31.52 12.98 31.62 13.08 ;
        RECT 31.52 12.74 31.62 12.84 ;
        RECT 31.52 12.5 31.62 12.6 ;
        RECT 31.52 12.26 31.62 12.36 ;
        RECT 31.52 12.02 31.62 12.12 ;
        RECT 31.72 13.7 31.82 13.8 ;
        RECT 31.72 13.46 31.82 13.56 ;
        RECT 31.72 13.22 31.82 13.32 ;
        RECT 31.72 12.98 31.82 13.08 ;
        RECT 31.72 12.74 31.82 12.84 ;
        RECT 31.72 12.5 31.82 12.6 ;
        RECT 31.72 12.26 31.82 12.36 ;
        RECT 31.72 12.02 31.82 12.12 ;
        RECT 31.92 13.7 32.02 13.8 ;
        RECT 31.92 13.46 32.02 13.56 ;
        RECT 31.92 13.22 32.02 13.32 ;
        RECT 31.92 12.98 32.02 13.08 ;
        RECT 31.92 12.74 32.02 12.84 ;
        RECT 31.92 12.5 32.02 12.6 ;
        RECT 31.92 12.26 32.02 12.36 ;
        RECT 31.92 12.02 32.02 12.12 ;
        RECT 32.12 13.7 32.22 13.8 ;
        RECT 32.12 13.46 32.22 13.56 ;
        RECT 32.12 13.22 32.22 13.32 ;
        RECT 32.12 12.98 32.22 13.08 ;
        RECT 32.12 12.74 32.22 12.84 ;
        RECT 32.12 12.5 32.22 12.6 ;
        RECT 32.12 12.26 32.22 12.36 ;
        RECT 32.12 12.02 32.22 12.12 ;
        RECT 32.32 13.7 32.42 13.8 ;
        RECT 32.32 13.46 32.42 13.56 ;
        RECT 32.32 13.22 32.42 13.32 ;
        RECT 32.32 12.98 32.42 13.08 ;
        RECT 32.32 12.74 32.42 12.84 ;
        RECT 32.32 12.5 32.42 12.6 ;
        RECT 32.32 12.26 32.42 12.36 ;
        RECT 32.32 12.02 32.42 12.12 ;
        RECT 32.52 13.7 32.62 13.8 ;
        RECT 32.52 13.46 32.62 13.56 ;
        RECT 32.52 13.22 32.62 13.32 ;
        RECT 32.52 12.98 32.62 13.08 ;
        RECT 32.52 12.74 32.62 12.84 ;
        RECT 32.52 12.5 32.62 12.6 ;
        RECT 32.52 12.26 32.62 12.36 ;
        RECT 32.52 12.02 32.62 12.12 ;
    END
    PORT
      LAYER M1 ;
        RECT -25 43.37 -20 48.375 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.77 43.515 33.66 44.415 ;
      LAYER M1 ;
        RECT 29.98 43.37 34.97 48.37 ;
      LAYER M2 ;
        RECT 32.77 43.515 33.66 44.415 ;
      LAYER VIA1 ;
        RECT 29.92 44.275 30.02 44.375 ;
        RECT 29.92 44.035 30.02 44.135 ;
        RECT 29.92 43.795 30.02 43.895 ;
        RECT 29.92 43.555 30.02 43.655 ;
        RECT 30.12 44.275 30.22 44.375 ;
        RECT 30.12 44.035 30.22 44.135 ;
        RECT 30.12 43.795 30.22 43.895 ;
        RECT 30.12 43.555 30.22 43.655 ;
        RECT 30.32 44.275 30.42 44.375 ;
        RECT 30.32 44.035 30.42 44.135 ;
        RECT 30.32 43.795 30.42 43.895 ;
        RECT 30.32 43.555 30.42 43.655 ;
        RECT 30.52 44.275 30.62 44.375 ;
        RECT 30.52 44.035 30.62 44.135 ;
        RECT 30.52 43.795 30.62 43.895 ;
        RECT 30.52 43.555 30.62 43.655 ;
        RECT 30.72 44.275 30.82 44.375 ;
        RECT 30.72 44.035 30.82 44.135 ;
        RECT 30.72 43.795 30.82 43.895 ;
        RECT 30.72 43.555 30.82 43.655 ;
        RECT 30.92 44.275 31.02 44.375 ;
        RECT 30.92 44.035 31.02 44.135 ;
        RECT 30.92 43.795 31.02 43.895 ;
        RECT 30.92 43.555 31.02 43.655 ;
        RECT 31.12 44.275 31.22 44.375 ;
        RECT 31.12 44.035 31.22 44.135 ;
        RECT 31.12 43.795 31.22 43.895 ;
        RECT 31.12 43.555 31.22 43.655 ;
        RECT 31.32 44.275 31.42 44.375 ;
        RECT 31.32 44.035 31.42 44.135 ;
        RECT 31.32 43.795 31.42 43.895 ;
        RECT 31.32 43.555 31.42 43.655 ;
        RECT 31.52 44.275 31.62 44.375 ;
        RECT 31.52 44.035 31.62 44.135 ;
        RECT 31.52 43.795 31.62 43.895 ;
        RECT 31.52 43.555 31.62 43.655 ;
        RECT 31.72 44.275 31.82 44.375 ;
        RECT 31.72 44.035 31.82 44.135 ;
        RECT 31.72 43.795 31.82 43.895 ;
        RECT 31.72 43.555 31.82 43.655 ;
        RECT 31.92 44.275 32.02 44.375 ;
        RECT 31.92 44.035 32.02 44.135 ;
        RECT 31.92 43.795 32.02 43.895 ;
        RECT 31.92 43.555 32.02 43.655 ;
        RECT 32.12 44.275 32.22 44.375 ;
        RECT 32.12 44.035 32.22 44.135 ;
        RECT 32.12 43.795 32.22 43.895 ;
        RECT 32.12 43.555 32.22 43.655 ;
        RECT 32.32 44.275 32.42 44.375 ;
        RECT 32.32 44.035 32.42 44.135 ;
        RECT 32.32 43.795 32.42 43.895 ;
        RECT 32.32 43.555 32.42 43.655 ;
        RECT 32.52 44.275 32.62 44.375 ;
        RECT 32.52 44.035 32.62 44.135 ;
        RECT 32.52 43.795 32.62 43.895 ;
        RECT 32.52 43.555 32.62 43.655 ;
        RECT 32.72 44.275 32.82 44.375 ;
        RECT 32.72 44.035 32.82 44.135 ;
        RECT 32.72 43.795 32.82 43.895 ;
        RECT 32.72 43.555 32.82 43.655 ;
        RECT 32.92 44.275 33.02 44.375 ;
        RECT 32.92 44.035 33.02 44.135 ;
        RECT 32.92 43.795 33.02 43.895 ;
        RECT 32.92 43.555 33.02 43.655 ;
        RECT 33.12 44.275 33.22 44.375 ;
        RECT 33.12 44.035 33.22 44.135 ;
        RECT 33.12 43.795 33.22 43.895 ;
        RECT 33.12 43.555 33.22 43.655 ;
        RECT 33.32 44.275 33.42 44.375 ;
        RECT 33.32 44.035 33.42 44.135 ;
        RECT 33.32 43.795 33.42 43.895 ;
        RECT 33.32 43.555 33.42 43.655 ;
        RECT 33.52 44.275 33.62 44.375 ;
        RECT 33.52 44.035 33.62 44.135 ;
        RECT 33.52 43.795 33.62 43.895 ;
        RECT 33.52 43.555 33.62 43.655 ;
      LAYER VIA2 ;
        RECT 29.92 44.275 30.02 44.375 ;
        RECT 29.92 44.035 30.02 44.135 ;
        RECT 29.92 43.795 30.02 43.895 ;
        RECT 29.92 43.555 30.02 43.655 ;
        RECT 30.12 44.275 30.22 44.375 ;
        RECT 30.12 44.035 30.22 44.135 ;
        RECT 30.12 43.795 30.22 43.895 ;
        RECT 30.12 43.555 30.22 43.655 ;
        RECT 30.32 44.275 30.42 44.375 ;
        RECT 30.32 44.035 30.42 44.135 ;
        RECT 30.32 43.795 30.42 43.895 ;
        RECT 30.32 43.555 30.42 43.655 ;
        RECT 30.52 44.275 30.62 44.375 ;
        RECT 30.52 44.035 30.62 44.135 ;
        RECT 30.52 43.795 30.62 43.895 ;
        RECT 30.52 43.555 30.62 43.655 ;
        RECT 30.72 44.275 30.82 44.375 ;
        RECT 30.72 44.035 30.82 44.135 ;
        RECT 30.72 43.795 30.82 43.895 ;
        RECT 30.72 43.555 30.82 43.655 ;
        RECT 30.92 44.275 31.02 44.375 ;
        RECT 30.92 44.035 31.02 44.135 ;
        RECT 30.92 43.795 31.02 43.895 ;
        RECT 30.92 43.555 31.02 43.655 ;
        RECT 31.12 44.275 31.22 44.375 ;
        RECT 31.12 44.035 31.22 44.135 ;
        RECT 31.12 43.795 31.22 43.895 ;
        RECT 31.12 43.555 31.22 43.655 ;
        RECT 31.32 44.275 31.42 44.375 ;
        RECT 31.32 44.035 31.42 44.135 ;
        RECT 31.32 43.795 31.42 43.895 ;
        RECT 31.32 43.555 31.42 43.655 ;
        RECT 31.52 44.275 31.62 44.375 ;
        RECT 31.52 44.035 31.62 44.135 ;
        RECT 31.52 43.795 31.62 43.895 ;
        RECT 31.52 43.555 31.62 43.655 ;
        RECT 31.72 44.275 31.82 44.375 ;
        RECT 31.72 44.035 31.82 44.135 ;
        RECT 31.72 43.795 31.82 43.895 ;
        RECT 31.72 43.555 31.82 43.655 ;
        RECT 31.92 44.275 32.02 44.375 ;
        RECT 31.92 44.035 32.02 44.135 ;
        RECT 31.92 43.795 32.02 43.895 ;
        RECT 31.92 43.555 32.02 43.655 ;
        RECT 32.12 44.275 32.22 44.375 ;
        RECT 32.12 44.035 32.22 44.135 ;
        RECT 32.12 43.795 32.22 43.895 ;
        RECT 32.12 43.555 32.22 43.655 ;
        RECT 32.32 44.275 32.42 44.375 ;
        RECT 32.32 44.035 32.42 44.135 ;
        RECT 32.32 43.795 32.42 43.895 ;
        RECT 32.32 43.555 32.42 43.655 ;
        RECT 32.52 44.275 32.62 44.375 ;
        RECT 32.52 44.035 32.62 44.135 ;
        RECT 32.52 43.795 32.62 43.895 ;
        RECT 32.52 43.555 32.62 43.655 ;
        RECT 32.72 44.275 32.82 44.375 ;
        RECT 32.72 44.035 32.82 44.135 ;
        RECT 32.72 43.795 32.82 43.895 ;
        RECT 32.72 43.555 32.82 43.655 ;
        RECT 32.92 44.275 33.02 44.375 ;
        RECT 32.92 44.035 33.02 44.135 ;
        RECT 32.92 43.795 33.02 43.895 ;
        RECT 32.92 43.555 33.02 43.655 ;
        RECT 33.12 44.275 33.22 44.375 ;
        RECT 33.12 44.035 33.22 44.135 ;
        RECT 33.12 43.795 33.22 43.895 ;
        RECT 33.12 43.555 33.22 43.655 ;
        RECT 33.32 44.275 33.42 44.375 ;
        RECT 33.32 44.035 33.42 44.135 ;
        RECT 33.32 43.795 33.42 43.895 ;
        RECT 33.32 43.555 33.42 43.655 ;
        RECT 33.52 44.275 33.62 44.375 ;
        RECT 33.52 44.035 33.62 44.135 ;
        RECT 33.52 43.795 33.62 43.895 ;
        RECT 33.52 43.555 33.62 43.655 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M1 ;
        RECT -20.51 14.515 -20.24 14.795 ;
    END
    PORT
      LAYER M1 ;
        RECT -20.51 2.545 -20.24 2.825 ;
    END
    PORT
      LAYER M1 ;
        RECT -25.03 -16.63 -20.04 -11.63 ;
    END
    PORT
      LAYER M1 ;
        RECT 29.98 -16.63 34.97 -11.63 ;
    END
    PORT
      LAYER M5 ;
        RECT 13 -12.88 14.38 -11.51 ;
      LAYER M4 ;
        RECT 13 -12.88 14.38 -12.19 ;
      LAYER M3 ;
        RECT 13 -12.88 14.38 -12.19 ;
      LAYER M2 ;
        RECT 13 -12.88 14.38 -12.19 ;
      LAYER VIA1 ;
        RECT 13.04 -11.84 13.14 -11.74 ;
        RECT 13.04 -12.04 13.14 -11.94 ;
        RECT 13.04 -12.24 13.14 -12.14 ;
        RECT 13.04 -12.44 13.14 -12.34 ;
        RECT 13.04 -12.64 13.14 -12.54 ;
        RECT 13.04 -12.84 13.14 -12.74 ;
        RECT 13.28 -11.84 13.38 -11.74 ;
        RECT 13.28 -12.04 13.38 -11.94 ;
        RECT 13.28 -12.24 13.38 -12.14 ;
        RECT 13.28 -12.44 13.38 -12.34 ;
        RECT 13.28 -12.64 13.38 -12.54 ;
        RECT 13.28 -12.84 13.38 -12.74 ;
        RECT 13.52 -11.84 13.62 -11.74 ;
        RECT 13.52 -12.04 13.62 -11.94 ;
        RECT 13.52 -12.24 13.62 -12.14 ;
        RECT 13.52 -12.44 13.62 -12.34 ;
        RECT 13.52 -12.64 13.62 -12.54 ;
        RECT 13.52 -12.84 13.62 -12.74 ;
        RECT 13.76 -11.84 13.86 -11.74 ;
        RECT 13.76 -12.04 13.86 -11.94 ;
        RECT 13.76 -12.24 13.86 -12.14 ;
        RECT 13.76 -12.44 13.86 -12.34 ;
        RECT 13.76 -12.64 13.86 -12.54 ;
        RECT 13.76 -12.84 13.86 -12.74 ;
        RECT 14 -11.84 14.1 -11.74 ;
        RECT 14 -12.04 14.1 -11.94 ;
        RECT 14 -12.24 14.1 -12.14 ;
        RECT 14 -12.44 14.1 -12.34 ;
        RECT 14 -12.64 14.1 -12.54 ;
        RECT 14 -12.84 14.1 -12.74 ;
        RECT 14.24 -11.84 14.34 -11.74 ;
        RECT 14.24 -12.04 14.34 -11.94 ;
        RECT 14.24 -12.24 14.34 -12.14 ;
        RECT 14.24 -12.44 14.34 -12.34 ;
        RECT 14.24 -12.64 14.34 -12.54 ;
        RECT 14.24 -12.84 14.34 -12.74 ;
      LAYER VIA2 ;
        RECT 13.04 -11.84 13.14 -11.74 ;
        RECT 13.04 -12.04 13.14 -11.94 ;
        RECT 13.04 -12.24 13.14 -12.14 ;
        RECT 13.04 -12.44 13.14 -12.34 ;
        RECT 13.04 -12.64 13.14 -12.54 ;
        RECT 13.04 -12.84 13.14 -12.74 ;
        RECT 13.28 -11.84 13.38 -11.74 ;
        RECT 13.28 -12.04 13.38 -11.94 ;
        RECT 13.28 -12.24 13.38 -12.14 ;
        RECT 13.28 -12.44 13.38 -12.34 ;
        RECT 13.28 -12.64 13.38 -12.54 ;
        RECT 13.28 -12.84 13.38 -12.74 ;
        RECT 13.52 -11.84 13.62 -11.74 ;
        RECT 13.52 -12.04 13.62 -11.94 ;
        RECT 13.52 -12.24 13.62 -12.14 ;
        RECT 13.52 -12.44 13.62 -12.34 ;
        RECT 13.52 -12.64 13.62 -12.54 ;
        RECT 13.52 -12.84 13.62 -12.74 ;
        RECT 13.76 -11.84 13.86 -11.74 ;
        RECT 13.76 -12.04 13.86 -11.94 ;
        RECT 13.76 -12.24 13.86 -12.14 ;
        RECT 13.76 -12.44 13.86 -12.34 ;
        RECT 13.76 -12.64 13.86 -12.54 ;
        RECT 13.76 -12.84 13.86 -12.74 ;
        RECT 14 -11.84 14.1 -11.74 ;
        RECT 14 -12.04 14.1 -11.94 ;
        RECT 14 -12.24 14.1 -12.14 ;
        RECT 14 -12.44 14.1 -12.34 ;
        RECT 14 -12.64 14.1 -12.54 ;
        RECT 14 -12.84 14.1 -12.74 ;
        RECT 14.24 -11.84 14.34 -11.74 ;
        RECT 14.24 -12.04 14.34 -11.94 ;
        RECT 14.24 -12.24 14.34 -12.14 ;
        RECT 14.24 -12.44 14.34 -12.34 ;
        RECT 14.24 -12.64 14.34 -12.54 ;
        RECT 14.24 -12.84 14.34 -12.74 ;
      LAYER VIA3 ;
        RECT 13.04 -11.84 13.14 -11.74 ;
        RECT 13.04 -12.04 13.14 -11.94 ;
        RECT 13.04 -12.24 13.14 -12.14 ;
        RECT 13.04 -12.44 13.14 -12.34 ;
        RECT 13.04 -12.64 13.14 -12.54 ;
        RECT 13.04 -12.84 13.14 -12.74 ;
        RECT 13.28 -11.84 13.38 -11.74 ;
        RECT 13.28 -12.04 13.38 -11.94 ;
        RECT 13.28 -12.24 13.38 -12.14 ;
        RECT 13.28 -12.44 13.38 -12.34 ;
        RECT 13.28 -12.64 13.38 -12.54 ;
        RECT 13.28 -12.84 13.38 -12.74 ;
        RECT 13.52 -11.84 13.62 -11.74 ;
        RECT 13.52 -12.04 13.62 -11.94 ;
        RECT 13.52 -12.24 13.62 -12.14 ;
        RECT 13.52 -12.44 13.62 -12.34 ;
        RECT 13.52 -12.64 13.62 -12.54 ;
        RECT 13.52 -12.84 13.62 -12.74 ;
        RECT 13.76 -11.84 13.86 -11.74 ;
        RECT 13.76 -12.04 13.86 -11.94 ;
        RECT 13.76 -12.24 13.86 -12.14 ;
        RECT 13.76 -12.44 13.86 -12.34 ;
        RECT 13.76 -12.64 13.86 -12.54 ;
        RECT 13.76 -12.84 13.86 -12.74 ;
        RECT 14 -11.84 14.1 -11.74 ;
        RECT 14 -12.04 14.1 -11.94 ;
        RECT 14 -12.24 14.1 -12.14 ;
        RECT 14 -12.44 14.1 -12.34 ;
        RECT 14 -12.64 14.1 -12.54 ;
        RECT 14 -12.84 14.1 -12.74 ;
        RECT 14.24 -11.84 14.34 -11.74 ;
        RECT 14.24 -12.04 14.34 -11.94 ;
        RECT 14.24 -12.24 14.34 -12.14 ;
        RECT 14.24 -12.44 14.34 -12.34 ;
        RECT 14.24 -12.64 14.34 -12.54 ;
        RECT 14.24 -12.84 14.34 -12.74 ;
      LAYER VIA4 ;
        RECT 13.04 -11.84 13.14 -11.74 ;
        RECT 13.04 -12.04 13.14 -11.94 ;
        RECT 13.04 -12.24 13.14 -12.14 ;
        RECT 13.04 -12.44 13.14 -12.34 ;
        RECT 13.04 -12.64 13.14 -12.54 ;
        RECT 13.04 -12.84 13.14 -12.74 ;
        RECT 13.28 -11.84 13.38 -11.74 ;
        RECT 13.28 -12.04 13.38 -11.94 ;
        RECT 13.28 -12.24 13.38 -12.14 ;
        RECT 13.28 -12.44 13.38 -12.34 ;
        RECT 13.28 -12.64 13.38 -12.54 ;
        RECT 13.28 -12.84 13.38 -12.74 ;
        RECT 13.52 -11.84 13.62 -11.74 ;
        RECT 13.52 -12.04 13.62 -11.94 ;
        RECT 13.52 -12.24 13.62 -12.14 ;
        RECT 13.52 -12.44 13.62 -12.34 ;
        RECT 13.52 -12.64 13.62 -12.54 ;
        RECT 13.52 -12.84 13.62 -12.74 ;
        RECT 13.76 -11.84 13.86 -11.74 ;
        RECT 13.76 -12.04 13.86 -11.94 ;
        RECT 13.76 -12.24 13.86 -12.14 ;
        RECT 13.76 -12.44 13.86 -12.34 ;
        RECT 13.76 -12.64 13.86 -12.54 ;
        RECT 13.76 -12.84 13.86 -12.74 ;
        RECT 14 -11.84 14.1 -11.74 ;
        RECT 14 -12.04 14.1 -11.94 ;
        RECT 14 -12.24 14.1 -12.14 ;
        RECT 14 -12.44 14.1 -12.34 ;
        RECT 14 -12.64 14.1 -12.54 ;
        RECT 14 -12.84 14.1 -12.74 ;
        RECT 14.24 -11.84 14.34 -11.74 ;
        RECT 14.24 -12.04 14.34 -11.94 ;
        RECT 14.24 -12.24 14.34 -12.14 ;
        RECT 14.24 -12.44 14.34 -12.34 ;
        RECT 14.24 -12.64 14.34 -12.54 ;
        RECT 14.24 -12.84 14.34 -12.74 ;
    END
  END GND
  PIN VOUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 17.4436 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 170.9008 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 136422 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30624 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1975680 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA5 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA6 ;
    ANTENNAPARTIALCUTAREA 1.0368 LAYER VIA7 ;
    PORT
      LAYER M2 ;
        RECT 33.225 9.435 34.365 10.575 ;
    END
  END VOUT
  PIN VINm
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2698 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 1.74935 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 56276 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 45430 LAYER M2 ;
    ANTENNAPARTIALCUTAREA 0.03 LAYER VIA2 ;
    PORT
      LAYER M2 ;
        RECT -23.575 7.085 -23.395 7.265 ;
    END
  END VINm
  PIN VINp
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.008 LAYER M3 ;
    ANTENNAPARTIALMETALAREA 10.9668 LAYER M2 ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M4 ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M5 ;
    ANTENNAPARTIALMETALAREA 1.7328 LAYER M6 ;
    ANTENNAPARTIALMETALAREA 2.5376 LAYER M7 ;
    ANTENNAPARTIALMETALAREA 86.8384 LAYER M8 ;
    ANTENNAPARTIALMETALSIDEAREA 83160 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 251680 LAYER M2 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M5 ;
    ANTENNAPARTIALMETALSIDEAREA 26752 LAYER M6 ;
    ANTENNAPARTIALMETALSIDEAREA 30624 LAYER M7 ;
    ANTENNAPARTIALMETALSIDEAREA 1064160 LAYER M8 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA3 ;
    ANTENNAPARTIALCUTAREA 0.43 LAYER VIA2 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA4 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA5 ;
    ANTENNAPARTIALCUTAREA 0.4 LAYER VIA6 ;
    ANTENNAPARTIALCUTAREA 1.0368 LAYER VIA7 ;
    PORT
      LAYER M2 ;
        RECT -23.575 5.95 -23.395 6.13 ;
    END
  END VINp
  OBS
    LAYER M1 ;
      RECT -22.71 37.985 33.81 38.845 ;
      RECT 32.95 -10.13 33.81 38.845 ;
      RECT 24.64 31.87 25.64 38.845 ;
      RECT 13.48 37.665 14.86 38.845 ;
      RECT -20.395 34.855 3.695 38.845 ;
      RECT -22.71 -10.13 -21.85 38.845 ;
      RECT 24.64 31.87 28.85 32.87 ;
      RECT 28.64 30.49 28.85 32.87 ;
      RECT 27.89 30.49 28.08 32.87 ;
      RECT 27.27 30.49 27.46 32.87 ;
      RECT 26.65 30.49 26.84 32.87 ;
      RECT 26.03 30.49 26.22 32.87 ;
      RECT 25.41 30.49 25.6 38.845 ;
      RECT 24.64 30.49 24.85 38.845 ;
      RECT -22.71 -9.56 -19.78 -0.42 ;
      RECT 21.285 7.825 23.525 16.965 ;
      RECT 2.99 16.135 4.91 16.305 ;
      RECT 4.74 8.265 4.91 16.305 ;
      RECT 2.99 8.265 3.16 16.305 ;
      RECT -8.205 14.02 -6.285 14.19 ;
      RECT -6.455 6.66 -6.285 14.19 ;
      RECT -8.205 6.66 -8.035 14.19 ;
      RECT 4.74 12.585 23.525 13.085 ;
      RECT 3.4 8.935 4.5 9.275 ;
      RECT 3.825 4.985 4.075 9.275 ;
      RECT 2.99 8.265 4.91 8.435 ;
      RECT -17.66 6.54 -9.54 8.32 ;
      RECT -10.04 -0.92 -9.54 8.32 ;
      RECT -7.795 7.14 -6.695 7.49 ;
      RECT -7.37 4.985 -7.12 7.49 ;
      RECT -8.205 6.66 -6.285 6.83 ;
      RECT -16.945 5.33 -11.095 5.54 ;
      RECT -11.305 -0.12 -11.095 5.54 ;
      RECT -14.125 3.28 -13.915 5.54 ;
      RECT -16.945 -0.12 -16.735 5.54 ;
      RECT -7.37 4.985 4.075 5.235 ;
      RECT -1.455 -16.63 -0.955 5.235 ;
      RECT -1.895 2.27 3.795 4.28 ;
      RECT -7.355 3.69 -3.045 3.86 ;
      RECT -3.215 -2.23 -3.045 3.86 ;
      RECT -4.825 2.2 -4.615 3.86 ;
      RECT -5.785 2.2 -5.575 3.86 ;
      RECT -7.355 -2.23 -7.185 3.86 ;
      RECT -10.04 -0.92 -8.26 3.16 ;
      RECT -1.895 -2.1 -0.575 4.28 ;
      RECT -14.125 -0.12 -13.915 2.14 ;
      RECT 0.12 1.21 3.81 1.38 ;
      RECT 3.64 -3.45 3.81 1.38 ;
      RECT 1.86 -0.17 2.07 1.38 ;
      RECT 0.12 -3.45 0.29 1.38 ;
      RECT -19.065 -0.12 -18.785 1.045 ;
      RECT -19.065 -0.12 -16.735 0.16 ;
      RECT -19.065 -0.12 -11.095 0.09 ;
      RECT -15.67 -2.07 -15.17 0.09 ;
      RECT -18.95 -1.25 -15.17 -0.75 ;
      RECT -9.26 -16.63 -8.76 3.16 ;
      RECT -18.95 -10.13 -18.45 -0.75 ;
      RECT -18.54 -16.63 -18.45 -0.75 ;
      RECT -17.705 -1.85 -10.375 -1.68 ;
      RECT -10.545 -8.47 -10.375 -1.68 ;
      RECT -13.395 -4.45 -13.185 -1.68 ;
      RECT -17.705 -8.47 -17.535 -1.68 ;
      RECT -16.725 -2.07 -14.115 -1.98 ;
      RECT -7.355 -2.23 -3.045 -2.06 ;
      RECT -14.27 -4.45 -14.05 -2.07 ;
      RECT -16.79 -4.45 -16.57 -2.07 ;
      RECT -15.11 -4.45 -14.89 -1.98 ;
      RECT -15.95 -4.45 -15.73 -1.98 ;
      RECT -6.185 -3.4 -5.685 -2.06 ;
      RECT -9.26 -2.985 -5.685 -2.485 ;
      RECT -7.8 -3.4 -2.24 -3.23 ;
      RECT -2.41 -9.36 -2.24 -3.23 ;
      RECT 0.12 -3.45 3.81 -3.28 ;
      RECT -4.33 -5.89 -4.12 -3.23 ;
      RECT -6.06 -3.73 -5.81 -2.06 ;
      RECT -7.8 -9.36 -7.63 -3.23 ;
      RECT 1.715 -5 2.215 -3.28 ;
      RECT -6.82 -3.73 -5.05 -3.64 ;
      RECT -5.14 -5.89 -5.05 -3.64 ;
      RECT -5.98 -5.89 -5.89 -2.06 ;
      RECT -6.82 -5.89 -6.73 -3.64 ;
      RECT 1.715 -4.375 4.625 -3.875 ;
      RECT 4.125 -16.63 4.625 -3.875 ;
      RECT -11.025 -6.225 -10.935 -4.355 ;
      RECT -11.865 -8.47 -11.775 -4.355 ;
      RECT -12.705 -6.225 -12.615 -4.355 ;
      RECT 0.07 -5 3.86 -4.83 ;
      RECT 3.69 -9.36 3.86 -4.83 ;
      RECT 2.71 -5.33 2.96 -4.83 ;
      RECT 1.86 -6.69 2.07 -3.28 ;
      RECT 0.97 -5.33 1.22 -4.83 ;
      RECT 0.07 -9.36 0.24 -4.83 ;
      RECT 2.37 -5.33 3.3 -5.24 ;
      RECT 3.21 -6.69 3.3 -5.24 ;
      RECT 0.63 -5.33 1.56 -5.24 ;
      RECT 1.47 -6.69 1.56 -5.24 ;
      RECT 2.37 -6.69 2.46 -5.24 ;
      RECT 0.63 -6.69 0.72 -5.24 ;
      RECT -13.395 -8.47 -13.185 -5.7 ;
      RECT -14.27 -8.08 -14.05 -5.7 ;
      RECT -15.11 -8.17 -14.89 -5.7 ;
      RECT -15.95 -8.17 -15.73 -5.7 ;
      RECT -16.79 -8.08 -16.57 -5.7 ;
      RECT -2.89 -6.925 -2.8 -5.875 ;
      RECT -3.73 -6.925 -3.64 -5.875 ;
      RECT -12.705 -6.225 -10.935 -6.135 ;
      RECT -11.94 -8.47 -11.69 -6.135 ;
      RECT -4.33 -9.36 -4.12 -6.7 ;
      RECT -5.14 -8.95 -5.05 -6.7 ;
      RECT -5.98 -9.36 -5.89 -6.7 ;
      RECT -6.82 -8.95 -6.73 -6.7 ;
      RECT 28.64 -9.095 28.85 -6.715 ;
      RECT 27.89 -9.095 28.08 -6.715 ;
      RECT 27.27 -9.095 27.46 -6.715 ;
      RECT 26.65 -9.095 26.84 -6.715 ;
      RECT 26.03 -9.095 26.22 -6.715 ;
      RECT 25.41 -16.63 25.6 -6.715 ;
      RECT 24.64 -16.63 24.85 -6.715 ;
      RECT -3.73 -6.925 -2.8 -6.835 ;
      RECT -3.385 -9.36 -3.135 -6.835 ;
      RECT 3.21 -8.95 3.3 -7.5 ;
      RECT 2.37 -8.95 2.46 -7.5 ;
      RECT 1.86 -16.63 2.07 -7.5 ;
      RECT 1.47 -8.95 1.56 -7.5 ;
      RECT 0.63 -8.95 0.72 -7.5 ;
      RECT -16.725 -8.17 -14.115 -8.08 ;
      RECT 24.64 -9.095 28.85 -8.095 ;
      RECT -15.67 -16.63 -15.17 -8.08 ;
      RECT -17.705 -8.47 -10.375 -8.3 ;
      RECT 2.37 -8.95 3.3 -8.86 ;
      RECT 0.63 -8.95 1.56 -8.86 ;
      RECT -6.82 -8.95 -5.05 -8.86 ;
      RECT 2.72 -9.36 2.97 -8.86 ;
      RECT 0.97 -9.36 1.22 -8.86 ;
      RECT -6.06 -9.36 -5.81 -8.86 ;
      RECT 24.64 -16.63 25.64 -8.095 ;
      RECT -14.43 -16.63 -9.89 -9.16 ;
      RECT 0.07 -9.36 3.86 -9.19 ;
      RECT -7.8 -9.36 -2.24 -9.19 ;
      RECT 1.715 -16.63 2.215 -9.19 ;
      RECT -5.5 -16.63 -5 -9.19 ;
      RECT -18.54 -16.63 28.48 -10.77 ;
      RECT -18.5 43.37 28.48 48.37 ;
      RECT -19.065 4.325 -18.785 13.015 ;
    LAYER M1 SPACING 0.09 ;
      RECT -19.82 -16.63 29.8 48.375 ;
      RECT -25.03 14.975 34.97 43.19 ;
      RECT -20.06 -11.45 34.97 43.19 ;
      RECT -20.46 14.94 -20.16 43.19 ;
      RECT -25.03 -11.45 -20.69 43.19 ;
      RECT -20.46 2.97 -20.16 14.37 ;
      RECT -25.03 3.005 34.97 14.335 ;
      RECT -20.46 -11.45 -20.16 2.4 ;
      RECT -25.03 -11.45 34.97 2.365 ;
      RECT -19.86 -16.63 29.8 43.19 ;
    LAYER M2 ;
      RECT 29.68 43.515 31.27 44.415 ;
    LAYER M2 SPACING 0.1 ;
      RECT -19.81 -12 29.79 48.375 ;
      RECT 14.57 -16.63 29.79 48.375 ;
      RECT -19.81 43.515 32.58 44.415 ;
      RECT -25.03 14.985 34.97 43.18 ;
      RECT 34.555 -11.44 34.97 43.18 ;
      RECT -20.4 14.95 34.97 43.18 ;
      RECT 32.85 10.765 34.97 43.18 ;
      RECT -25.03 7.455 -20.7 43.18 ;
      RECT -20.05 14.03 34.97 43.18 ;
      RECT -20.4 14.03 34.97 14.36 ;
      RECT -23.205 3.015 30.62 14.325 ;
      RECT -20.05 -11.44 33.035 11.79 ;
      RECT -20.05 -11.44 34.97 9.245 ;
      RECT -25.03 -11.44 -23.765 43.18 ;
      RECT -25.03 6.32 34.97 6.895 ;
      RECT -25.03 -11.44 -20.7 5.76 ;
      RECT -20.4 2.98 -20.22 14.36 ;
      RECT -20.4 -11.44 -20.22 2.39 ;
      RECT -25.03 -11.44 34.97 2.355 ;
      RECT -19.85 -16.63 12.81 43.18 ;
      RECT -19.85 -16.63 29.79 -13.07 ;
    LAYER M3 SPACING 0.1 ;
      RECT -25.03 44.605 34.97 48.375 ;
      RECT 34.555 -16.63 34.97 48.375 ;
      RECT 33.85 10.765 34.97 48.375 ;
      RECT -25.03 7.455 32.58 48.375 ;
      RECT -25.03 10.765 34.97 43.325 ;
      RECT -25.03 7.455 33.035 43.325 ;
      RECT 14.57 -16.63 34.97 9.245 ;
      RECT -23.205 -12 34.97 9.245 ;
      RECT -25.03 -16.63 -23.765 48.375 ;
      RECT -25.03 6.32 34.97 6.895 ;
      RECT -25.03 -16.63 12.81 5.76 ;
      RECT -25.03 -16.63 34.97 -13.07 ;
    LAYER M4 ;
      RECT 21.9 29.99 22.28 31.13 ;
      RECT 21.43 -4.37 21.81 -3.23 ;
      RECT 21 24.425 21.38 25.565 ;
      RECT 21 35.525 21.38 36.665 ;
      RECT 20.52 -9.925 20.9 -8.785 ;
      RECT 20.52 1.175 20.9 2.315 ;
      RECT 18.58 7.895 18.96 9.035 ;
      RECT 18.575 17.74 18.955 18.88 ;
      RECT 17.67 4.845 18.05 5.985 ;
      RECT 17.67 10.945 18.05 12.085 ;
      RECT 17.665 14.7 18.045 15.84 ;
      RECT 17.665 20.8 18.045 21.94 ;
      RECT 13.48 37.665 14.86 38.845 ;
      RECT 13 -11.94 14.38 -11.7 ;
    LAYER M5 ;
      RECT 13.48 21.65 14.86 38.845 ;
      RECT 7.905 36.375 20.425 36.805 ;
      RECT 17.165 33.545 18.365 36.805 ;
      RECT 15.365 31.745 16.565 36.805 ;
      RECT 11.765 31.745 12.965 36.805 ;
      RECT 9.965 33.545 11.165 36.805 ;
      RECT 17.165 33.545 20.425 34.745 ;
      RECT 7.905 33.545 11.165 34.745 ;
      RECT 15.365 31.745 20.425 32.945 ;
      RECT 7.905 31.745 12.965 32.945 ;
      RECT 7.905 29.945 20.425 31.145 ;
      RECT 15.365 28.145 20.425 29.345 ;
      RECT 7.905 28.145 12.965 29.345 ;
      RECT 11.765 24.285 12.965 29.345 ;
      RECT 15.365 24.285 16.565 29.345 ;
      RECT 17.165 26.345 20.425 27.545 ;
      RECT 7.905 26.345 11.165 27.545 ;
      RECT 9.965 24.285 11.165 27.545 ;
      RECT 17.165 24.285 18.365 27.545 ;
      RECT 7.905 24.285 20.425 24.715 ;
      RECT 9.575 21.65 17.095 22.08 ;
      RECT 14.535 19.52 15.735 22.08 ;
      RECT 12.735 14.56 13.935 22.08 ;
      RECT 10.935 19.52 12.135 22.08 ;
      RECT 14.535 19.52 17.095 20.72 ;
      RECT 9.575 19.52 12.135 20.72 ;
      RECT 9.575 17.72 17.095 18.92 ;
      RECT 14.535 15.92 17.095 17.12 ;
      RECT 9.575 15.92 12.135 17.12 ;
      RECT 10.935 14.56 12.135 17.12 ;
      RECT 14.535 14.56 15.735 17.12 ;
      RECT 9.575 14.56 17.095 14.99 ;
      RECT 9.58 11.795 17.1 12.225 ;
      RECT 14.54 9.665 15.74 12.225 ;
      RECT 12.74 4.705 13.94 12.225 ;
      RECT 10.94 9.665 12.14 12.225 ;
      RECT 14.54 9.665 17.1 10.865 ;
      RECT 9.58 9.665 12.14 10.865 ;
      RECT 9.58 7.865 17.1 9.065 ;
      RECT 14.54 6.065 17.1 7.265 ;
      RECT 9.58 6.065 12.14 7.265 ;
      RECT 10.94 4.705 12.14 7.265 ;
      RECT 14.54 4.705 15.74 7.265 ;
      RECT 9.58 4.705 17.1 5.135 ;
      RECT 13 -11.26 14.38 5.135 ;
      RECT 7.43 2.025 19.95 2.455 ;
      RECT 16.69 -0.805 17.89 2.455 ;
      RECT 14.89 -2.605 16.09 2.455 ;
      RECT 11.29 -2.605 12.49 2.455 ;
      RECT 9.49 -0.805 10.69 2.455 ;
      RECT 16.69 -0.805 19.95 0.395 ;
      RECT 7.43 -0.805 10.69 0.395 ;
      RECT 14.89 -2.605 19.95 -1.405 ;
      RECT 7.43 -2.605 12.49 -1.405 ;
      RECT 7.43 -4.405 19.95 -3.205 ;
      RECT 14.89 -6.205 19.95 -5.005 ;
      RECT 7.43 -6.205 12.49 -5.005 ;
      RECT 11.29 -10.065 12.49 -5.005 ;
      RECT 14.89 -10.065 16.09 -5.005 ;
      RECT 16.69 -8.005 19.95 -6.805 ;
      RECT 7.43 -8.005 10.69 -6.805 ;
      RECT 9.49 -10.065 10.69 -6.805 ;
      RECT 16.69 -10.065 17.89 -6.805 ;
      RECT 7.43 -10.065 19.95 -9.635 ;
      RECT 21.9 29.99 22.28 31.13 ;
      RECT 21.43 -4.37 21.81 -3.23 ;
      RECT 21 24.425 21.38 25.565 ;
      RECT 21 35.525 21.38 36.665 ;
      RECT 20.52 -9.925 20.9 -8.785 ;
      RECT 20.52 1.175 20.9 2.315 ;
      RECT 18.58 7.895 18.96 9.035 ;
      RECT 18.575 17.74 18.955 18.88 ;
      RECT 17.67 4.845 18.05 5.985 ;
      RECT 17.67 10.945 18.05 12.085 ;
      RECT 17.665 14.7 18.045 15.84 ;
      RECT 17.665 20.8 18.045 21.94 ;
    LAYER M6 ;
      RECT 14.465 29.045 20.425 30.245 ;
      RECT 7.905 29.045 13.865 30.245 ;
      RECT 12.665 24.285 13.865 30.245 ;
      RECT 14.465 24.285 15.665 30.245 ;
      RECT 16.265 27.245 20.425 28.445 ;
      RECT 7.905 27.245 12.065 28.445 ;
      RECT 10.865 24.285 12.065 28.445 ;
      RECT 16.265 24.285 17.465 28.445 ;
      RECT 18.065 24.285 20.425 26.645 ;
      RECT 7.905 24.285 10.265 26.645 ;
      RECT 7.905 24.285 20.425 24.715 ;
      RECT 7.905 36.375 20.425 36.805 ;
      RECT 18.065 34.445 20.425 36.805 ;
      RECT 16.265 32.645 17.465 36.805 ;
      RECT 14.465 30.845 15.665 36.805 ;
      RECT 12.665 30.845 13.865 36.805 ;
      RECT 10.865 32.645 12.065 36.805 ;
      RECT 7.905 34.445 10.265 36.805 ;
      RECT 16.265 32.645 20.425 33.845 ;
      RECT 7.905 32.645 12.065 33.845 ;
      RECT 14.465 30.845 20.425 32.045 ;
      RECT 7.905 30.845 13.865 32.045 ;
      RECT 13.99 -5.305 19.95 -4.105 ;
      RECT 7.43 -5.305 13.39 -4.105 ;
      RECT 12.19 -10.065 13.39 -4.105 ;
      RECT 13.99 -10.065 15.19 -4.105 ;
      RECT 15.79 -7.105 19.95 -5.905 ;
      RECT 7.43 -7.105 11.59 -5.905 ;
      RECT 10.39 -10.065 11.59 -5.905 ;
      RECT 15.79 -10.065 16.99 -5.905 ;
      RECT 17.59 -10.065 19.95 -7.705 ;
      RECT 7.43 -10.065 9.79 -7.705 ;
      RECT 7.43 -10.065 19.95 -9.635 ;
      RECT 7.43 2.025 19.95 2.455 ;
      RECT 17.59 0.095 19.95 2.455 ;
      RECT 15.79 -1.705 16.99 2.455 ;
      RECT 13.99 -3.505 15.19 2.455 ;
      RECT 12.19 -3.505 13.39 2.455 ;
      RECT 10.39 -1.705 11.59 2.455 ;
      RECT 7.43 0.095 9.79 2.455 ;
      RECT 15.79 -1.705 19.95 -0.505 ;
      RECT 7.43 -1.705 11.59 -0.505 ;
      RECT 13.99 -3.505 19.95 -2.305 ;
      RECT 7.43 -3.505 13.39 -2.305 ;
      RECT 13.64 6.965 17.1 8.165 ;
      RECT 9.58 6.965 13.04 8.165 ;
      RECT 11.84 4.705 13.04 8.165 ;
      RECT 13.64 4.705 14.84 8.165 ;
      RECT 15.44 4.705 17.1 6.365 ;
      RECT 9.58 4.705 11.24 6.365 ;
      RECT 9.58 4.705 17.1 5.135 ;
      RECT 9.58 11.795 17.1 12.225 ;
      RECT 15.44 10.565 17.1 12.225 ;
      RECT 13.64 8.765 14.84 12.225 ;
      RECT 11.84 8.765 13.04 12.225 ;
      RECT 9.58 10.565 11.24 12.225 ;
      RECT 13.64 8.765 17.1 9.965 ;
      RECT 9.58 8.765 13.04 9.965 ;
      RECT 13.635 16.82 17.095 18.02 ;
      RECT 9.575 16.82 13.035 18.02 ;
      RECT 11.835 14.56 13.035 18.02 ;
      RECT 13.635 14.56 14.835 18.02 ;
      RECT 15.435 14.56 17.095 16.22 ;
      RECT 9.575 14.56 11.235 16.22 ;
      RECT 9.575 14.56 17.095 14.99 ;
      RECT 9.575 21.65 17.095 22.08 ;
      RECT 15.435 20.42 17.095 22.08 ;
      RECT 13.635 18.62 14.835 22.08 ;
      RECT 11.835 18.62 13.035 22.08 ;
      RECT 9.575 20.42 11.235 22.08 ;
      RECT 13.635 18.62 17.095 19.82 ;
      RECT 9.575 18.62 13.035 19.82 ;
      RECT 21.9 29.99 22.28 31.13 ;
      RECT 21.43 -4.37 21.81 -3.23 ;
      RECT 21 24.425 21.38 25.565 ;
      RECT 21 35.525 21.38 36.665 ;
      RECT 20.52 -9.925 20.9 -8.785 ;
      RECT 20.52 1.175 20.9 2.315 ;
      RECT 18.58 7.895 18.96 9.035 ;
      RECT 18.575 17.74 18.955 18.88 ;
      RECT 17.67 4.845 18.05 5.985 ;
      RECT 17.67 10.945 18.05 12.085 ;
      RECT 17.665 14.7 18.045 15.84 ;
      RECT 17.665 20.8 18.045 21.94 ;
    LAYER M7 ;
      RECT 21.83 29.95 22.35 31.17 ;
      RECT 21.36 -4.41 21.88 -3.19 ;
      RECT 20.93 24.385 21.45 25.605 ;
      RECT 20.93 35.485 21.45 36.705 ;
      RECT 20.45 -9.965 20.97 -8.745 ;
      RECT 20.45 1.135 20.97 2.355 ;
      RECT 18.51 7.855 19.03 9.075 ;
      RECT 18.505 17.7 19.025 18.92 ;
      RECT 17.6 4.805 18.12 6.025 ;
      RECT 17.6 10.905 18.12 12.125 ;
      RECT 17.595 14.66 18.115 15.88 ;
      RECT 17.595 20.76 18.115 21.98 ;
    LAYER M8 ;
      RECT 16.185 26.785 17.925 34.305 ;
      RECT 13.295 26.785 15.035 34.305 ;
      RECT 10.405 26.785 12.145 34.305 ;
      RECT 7.905 29.365 22.925 31.725 ;
      RECT 15.71 -7.565 17.45 -0.045 ;
      RECT 12.82 -7.565 14.56 -0.045 ;
      RECT 9.93 -7.565 11.67 -0.045 ;
      RECT 7.43 -4.985 22.45 -2.625 ;
      RECT 5.405 35.385 21.545 36.805 ;
      RECT 5.405 35.145 20.425 36.805 ;
      RECT 18.765 32.565 20.425 36.805 ;
      RECT 7.905 32.565 9.565 36.805 ;
      RECT 5.405 24.285 7.065 36.805 ;
      RECT 18.765 24.285 20.425 28.525 ;
      RECT 7.905 24.285 9.565 28.525 ;
      RECT 5.405 24.285 20.425 25.945 ;
      RECT 5.405 24.285 21.545 25.705 ;
      RECT 4.93 1.035 21.07 2.455 ;
      RECT 4.93 0.795 19.95 2.455 ;
      RECT 18.29 -1.785 19.95 2.455 ;
      RECT 7.43 -1.785 9.09 2.455 ;
      RECT 4.93 -10.065 6.59 2.455 ;
      RECT 18.29 -10.065 19.95 -5.825 ;
      RECT 7.43 -10.065 9.09 -5.825 ;
      RECT 4.93 -10.065 19.95 -8.405 ;
      RECT 4.93 -10.065 21.07 -8.645 ;
      RECT 12.47 7.205 14.21 9.725 ;
      RECT 9.58 7.285 19.6 9.645 ;
      RECT 12.465 17.06 14.205 19.58 ;
      RECT 9.575 17.14 19.595 19.5 ;
      RECT 7.08 10.805 18.22 12.225 ;
      RECT 7.08 10.565 17.1 12.225 ;
      RECT 7.08 4.705 8.74 12.225 ;
      RECT 7.08 4.705 17.1 6.365 ;
      RECT 7.08 4.705 18.22 6.125 ;
      RECT 7.075 20.66 18.215 22.08 ;
      RECT 7.075 20.42 17.095 22.08 ;
      RECT 7.075 14.56 8.735 22.08 ;
      RECT 7.075 14.56 17.095 16.22 ;
      RECT 7.075 14.56 18.215 15.98 ;
  END
  PROPERTY pathCL "yes" ;
  PROPERTY arrayDisplay "Full" ;
  PROPERTY instLabel "master" ;
  PROPERTY startLevel 0 ;
  PROPERTY stopLevel 31 ;
  PROPERTY scrollPercent 25 ;
  PROPERTY gridSpacing 1 ;
  PROPERTY gridMultiple 5 ;
  PROPERTY xSnapSpacing 0.005 ;
  PROPERTY ySnapSpacing 0.005 ;
  PROPERTY snapMode "orthogonal" ;
  PROPERTY segSnapMode "orthogonal" ;
  PROPERTY instanceDrawingMode "BBox" ;
  PROPERTY lppVisibilityMode "donotCheckValidity" ;
  PROPERTY filterSize 6 ;
  PROPERTY filterSizeDrawingStyle "empty" ;
  PROPERTY displayResolution "Medium" ;
  PROPERTY dimmingScope "none" ;
  PROPERTY dimmingIntensity 50 ;
  PROPERTY autoZoomMode "Pan" ;
  PROPERTY autoZoomScale 90 ;
  PROPERTY mergeScope "pcells" ;
  PROPERTY viewNameList "spectre cmos_sch cmos.sch av_extracted schematic veriloga" ;
END X0814_opamp_N_P

END LIBRARY
